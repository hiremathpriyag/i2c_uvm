


   // dut wrapper including two interfaces 
     module dut_wrap();

    `include master_interface.sv
    `include slave_interface.sv

    endmodule

    

   
